library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
use ieee.std_logic_unsigned.all ;

entity mapp is
port (
x_now,y_now: in integer;
winn: in std_logic;
assign_mapwin:out std_logic;
assign_maze:out std_logic);
end mapp;
architecture lets_say of mapp is
type mazemap is array (0 to 119) of std_logic_vector(0 to 159);
constant the_map : mazemap := (
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000100000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000001000000000000000000100000000000000000000000000000000000010000",
"0011111111111111111111111000000000000000000100000000000000000100000000000000000001000000000000000001111111111111111111111111111111111111100000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000001111111111111111111111111111111111111100000000000000000001000000000000000011111111111111111111111111111111111111111111111111111111110000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000",
"0010000000000000000000001000000000000000000100000000000000000111111111111111111111111111111111111110000000000000000000111111111111111111100000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000",
"0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000110000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);

type bitwinmap is array (0 to 119) of std_logic_vector(0 to 159);
constant the_winmap : bitwinmap := (
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001100000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100001110000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100001111000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001111000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001111100000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111100000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001111110000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001111110000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001111111000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111111000000000000",
"0000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000",
"0000000000000000000000011111100000000011100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000110001111111100000000000",
"0000000000000000000011111000011111111100011000000000000000000000000000000000000000000000000000000000000000011111000000011100000000000000010110000000000000000000",
"0000000000000000001111000111100000000011100100000000000000000000000000000000000000000000000000000000000001111000111111100011000000000000010001111111100000000000",
"0000000000000000011100111000011111111100011010000000000000000000000000000000000000000000000000000000000011100111000000011100100000000000011110000000000000000000",
"0000000000000001111011000111100000000011100101000000000000000000000000000000000000000000000000000000000111011000111111100011011000000000011001111111110000000000",
"0000000000000011100100111000011111111100011010000000000000000000000000000000000000000000000000000000001110100111000000011100100100000000001010000000000000000000",
"0000000000000111011011000111100000000011100101100000000000000000000000000000000000000000000000000000011101011000111111100011011010000000001001111111110000000000",
"0000000000001110100100111000011111111100011010000000000000000000000001111111111000000000000000000000101010100111000000011100100101000000001110000000000000000000",
"0000000000011101011011000111100000000011100101100000000000000000001111100000000111000000000000000000110101011000111111100011011010000000001101111111111000000000",
"0000000000111010100100111000011111111100011010000000000000000000111100011111111000110000000000000001111010100111000000011100100101100000000100000000000000000000",
"0000000001110101011011000111100000000011100101000000000000000001110011100000000111001100000000000010100101011000111111100011011010010000000101111111111000000000",
"0000000010101010100100111000011111111100011010000000000000000111101100011111111000110010000000000010011010100111000000011100100101100000000110000000000000000000",
"0000000011010101011011000111100000000011100100000000000000001010010011100000000111001101000000000011100101011000110001100011011010011000000110111111111100000000",
"0000000101101010100100111000000000000000110000000000000000001101101100011111111000110010100000000101011010100111000000011100100101100000000010000000000000000000",
"0000000110010101011011000100000000000000000000000000000000011110010011100000000111001101010000000100100101011000000000001111011010011100000010111111111100000000",
"0000001011101010100100110000000000000000000000000000000000111001101100011111111000110010101000000101011010100100000000000110100101100000000011000000000000000000",
"0000001000010101011011000000000000000000000000000000000001010110010011100000000111001101010100000100100101011000000000000010011010011100000011011111111110000000",
"0000001111101010100100000000000000000000000000000000000001101001101100011111111000110010101000000101011010100100000000000011100101100010000001000000000000000000",
"0000010100010101011011000000000000000000000000000000000010110110010011100000000111001101010110000100100101011000000000000011011010011100000001011111111110000000",
"0000010011101010100100000000000000000000000000000000000010001001101100011111111000110010101000000101011010100100000000000001000101100010000001100000000000000000",
"0000010100010101011010000000000000000000000000000000000011110110010011100000001111001101010111000100100101011000000000000001011010011100000001101111111110000000",
"0000010011101010100100000000000000000000000000000000000101001001101100000000000110110010101000000101011010100100000000000001000101100010000000100000000001000000",
"0000010100010101011010000000000000000000000000000000000100110110010010000000000011001101010111100100100101011000000000000001011010011101000000101111111110000000",
"0000010011101010100100000000000000000000000000000000000101001001101100000000000001100010101000000111011010100100000000000001000101100010000000110000000001000000",
"0000010100010101011000000000000000000000000000000000000100110110010010000000000000101101010111100110100101011000000000000001011010011101000000110111111110100000",
"0000010011101010100100000000000000000000000000000000000101001001101100000000000000110010101000000010011010100110000000000001000101100010000000010000000001000000",
"0000010100010101011000000000000000000000000000000000000100110110010000000000000000110101010111110011100101011000000000000001011010011101000000010111111110100000",
"0000010011101010100100000000000000000000000000000000000101001001101100000000000000010010101000000011011010100111000000000001100101100010000000011000000001000000",
"0000010100010101011000000000000000000000000000000000000100110110010000000000000000010101010111110001100101011000100000000011111010011100000000011011111110100000",
"0000010011101010100110000000000000000000000000000000000101001001101110000000000000010010101000000001101010100111010000000111000101100010000000001000000001000000",
"0000010100010101011000000000000000000000000000000000000100110110010000000000000000010101010111110000110101011000101100011110111010011100000000001111111110100000",
"0000010011101010100110000000000000000000000000000000000111001001101110000000000000010010101000000000110010100111010011111001000101100000000000001100000001000000",
"0000010100010101011000000000000000000000000000000000000110110110010000000000000000010101010111110000011101011000101100000110111010011100000000000111111110100000",
"0000011011101010100110000000000000000000000000000000000010001001101111000000000000010010101000000000011010100111010011111001000101100000000000000110000001000000",
"0000011000010101011001000000000000000000000000000000000011110110010000000000000000011101010111110000001101011000101100000110111010011000000000000011111110000000",
"0000001011101010100110000000000000000000000000000000000011001001101111100000000000111010101000000000000110100111010011111001000101100000000000000001100000000000",
"0000001100010101011001000000000000000000000000000000000001110110010000010000000001110101010111110000000111011000101100000110111010010000000000000000011000000000",
"0000001101101010100110100000000000000000000000000000000001101001101111101000000011101010101000000000000011100111010011111001000101100000000000000000000000000000",
"0000000100010101011001000000000000000000000000000000000000110110010000010110000111010101010111100000000000111000101100000110111010000000000000000000000000000000",
"0000000111101010100110110000000000000000000000000000000000110001101111101001111110101010101000000000000000011111010011111001000100000000000000000000000000000000",
"0000000110010101011001000000000000000000000000000000000000011110010000010110000001010101010111000000000000001100101100000110111000000000000000000000000000000000",
"0000000010101010100110111000000000000000000000001111000000011001101111101001111110101010101000000000000000000011010011111001000000000000000000000000000000000000",
"0000000011010101011001000100000000000000000000111100110000001100010000010110000001010101010110000000000000000000011100000110000000000000000000000000000000000000",
"0000000011101010100110111010000000000000000001110011001000000111101111101001111110101010101000000000000000000000000000000000000000000000000000000000000000000000",
"0000000001100101011001000101000000000000000111101100110000000110010000010110000001010101010100000000000000000000000000000000000000000000000000000000000000000000",
"0000000000111010100110111010110000000000011110010011001100000011101111101001111110101010101000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000110101011001000101001110000011111001101100110000000001110000010110000001010101010000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000011010100110111010110001111111000110010011001100000000011111101001111110101010100000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000001101011001000101001110000000111001101100110000000000001100010110000001010101000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000001110100110111010110001111111000110010011001100000000000011101001111110101000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000111011001000101001110000000111001101100110000000000000000110110000001010000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000011100110111010110001111111000110010011001000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000001111001000101001110000000111001101100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000110110111010110001111111000110010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000011001000101001110000000111001101100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000001110111010110001111111000110010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000011000101001110000000111001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000111010110001111111000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000001101001110000000111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000011110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"

);
begin
process(x_now,y_now,winn)
begin
if (winn='0') then
	assign_mapwin<= '0';
	if y_now < 480 and x_now < 640 then
		assign_maze<= the_map(y_now/4)(x_now/4);
	else
		assign_maze<= '0';
	end if;

else 
	assign_maze<= '0';
	if y_now < 480 and x_now < 640 then
		assign_mapwin<= the_winmap(y_now/4)(x_now/4);
	else
		assign_mapwin<= '0';
	end if;
end if;
end process;

end lets_say;


LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all ;
USE ieee.std_logic_arith.all ;
USE ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity winning is
Port ( reset: in std_logic;
		 x_now,y_now : in integer;
		 assign: in std_logic;
		 win_res	: out std_logic;
		 win : out std_logic);
end winning ;

architecture Structural of winning is

signal gecici: std_logic:='0';
begin

process(x_now,y_now,assign,reset)
begin
if(reset='1') then 
gecici<='0';
win_res<='0';
elsif ((x_now<595 and x_now>=590) and (y_now<445 and y_now>=440)) then
win_res<='1';
 if(assign='1') then 
 gecici<='1';
 else
 gecici<='0';
 end if;
else 
gecici<=gecici;
win_res<='0';
end if;
end process;
win<=gecici;
end Structural;

LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all ;
USE ieee.std_logic_arith.all ;
USE ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity freq_div_2 is
Port ( clk : in std_logic;
slowed_clk : out std_logic);
end freq_div_2 ;

architecture Structural of freq_div_2 is

signal ara: std_logic_vector(1 downto 0);
signal not_ara: std_logic_vector(1 downto 0);
begin
not_ara(1)<= not ara(1);
not_ara(0)<= not ara(0);
u0: FDCE port map (C => clk, CE => '1', CLR => '0', D => not_ara(1), Q => ara(1));

u1: FDCE port map (C => ara(1), CE => '1', CLR => '0', D => not_ara(0), Q => ara(0));


slowed_clk <= ara(0);

end Structural;



LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all ;
USE ieee.std_logic_arith.all ;
USE ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity freq_div_20 is
Port ( clk : in std_logic;
slowed_clk : out std_logic);
end freq_div_20 ;

architecture Structural of freq_div_20 is

signal ara: std_logic_vector(19 downto 0);
signal not_ara: std_logic_vector(19 downto 0);
begin
not_ara(19)<= not ara(19);
not_ara(18)<= not ara(18);
not_ara(17)<= not ara(17);
not_ara(16)<= not ara(16);
not_ara(15)<= not ara(15);
not_ara(14)<= not ara(14);
not_ara(13)<= not ara(13);
not_ara(12)<= not ara(12);
not_ara(11)<= not ara(11);
not_ara(10)<= not ara(10);
not_ara(9)<= not ara(9);
not_ara(8)<= not ara(8);
not_ara(7)<= not ara(7);
not_ara(6)<= not ara(6);
not_ara(5)<= not ara(5);
not_ara(4)<= not ara(4);
not_ara(3)<= not ara(3);
not_ara(2)<= not ara(2);
not_ara(1)<= not ara(1);
not_ara(0)<= not ara(0);
u0: FDCE port map (C => clk, CE => '1', CLR => '0', D => not_ara(19), Q => ara(19));

c: for i in 1 to 19 generate
	u1to19: FDCE port map (C => ara(i), CE => '1', CLR => '0', D => not_ara(i-1), Q => ara(i-1));
end generate;

slowed_clk <= ara(0);

end Structural;

LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all ;
USE ieee.std_logic_arith.all ;
USE ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity shift_4 is
Port ( btn : in std_logic;
slowed_clk : in std_logic;
deb_out : out std_logic);
end shift_4 ;

architecture Structural of shift_4 is

signal ara : std_logic_vector (3 downto 0);

begin

s0: FDCE port map (C => slowed_clk, CE => '1', CLR => '0', D => btn, Q => ara(3));
s1: FDCE port map (C => slowed_clk, CE => '1', CLR => '0', D => ara(3), Q => ara(2));
s2: FDCE port map (C => slowed_clk, CE => '1', CLR => '0', D => ara(2), Q => ara(1));
s3: FDCE port map (C => slowed_clk, CE => '1', CLR => '0', D => ara(1), Q => ara(0));

deb_out <= ara(3) and ara(2) and ara(1) and ara(0);

end Structural;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


package square is 
procedure sq(signal x_now,y_now,xpos,ypos : IN INTEGER ;
signal assign : OUT std_logic );
end square;

package body square is 
procedure sq(signal x_now,y_now,xpos,ypos : IN INTEGER ;
signal assign : OUT std_logic )is
begin 
if( x_now>xpos and x_now<=(xpos+28) and y_now>ypos and y_now<=(ypos+28)) then
assign<='1';
else 
assign<='0';

end if;
end sq;
end square;




library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;
use IEEE.STD_LOGIC_ARITH.ALL;

entity vga2 is
    Port ( VL : in  STD_LOGIC;
           VU : in  STD_LOGIC;
           VD : in  STD_LOGIC;
			  VR : in  STD_LOGIC;
			  vclk : in  STD_LOGIC;
			  reset : in std_logic;
           vgahs,vgavs : out  STD_LOGIC;
           vgar : out  STD_LOGIC_vector(2 downto 0);
           vgag : out  STD_LOGIC_vector(2 downto 0);
           vgab : out  STD_LOGIC_vector(1 downto 0));
end vga2;

architecture Behavioral of vga2 is
use work.square.all;
signal slow,ssclk : std_logic;
signal dir : std_logic_vector(3 downto 0);
signal assign_sq,assign_mapwin,assign_maze,win_res,win : std_logic:='0';
signal hpos: integer range 0 to 799:=0;
signal vpos: integer range 0 to 520:=0;
signal refx:  INTEGER RANGE 0 to 799:=16;
signal refy : INTEGER RANGE 0 to 799:=16;
shared variable rgb : STD_LOGIC_VECTOR(7 downto 0):="11100000";


constant H_DISP : INTEGER :=640; 
constant H_FP	 :	INTEGER :=16;	
constant H_PW	 : INTEGER :=96;	
constant H_BP	 : INTEGER :=48;	


constant V_DISP : INTEGER :=480; 
constant V_FP	 :	INTEGER :=10;	
constant V_PW	 : INTEGER :=2;	
constant V_BP	 : INTEGER :=29;	


constant h_period : INTEGER := H_DISP + H_FP + H_PW + H_BP -1 ;
constant v_period : INTEGER := V_DISP + V_FP + V_PW + V_BP -1 ;

component winning 
Port ( reset: in std_logic;
		 x_now,y_now : in integer;
		 assign: in std_logic;
		 win_res	: out std_logic;
		 win : out std_logic);
end component ;

component mapp 
port (
x_now,y_now: in integer;
winn: in std_logic;
assign_mapwin:out std_logic;
assign_maze:out std_logic);
end component;

component freq_div_2 
Port ( clk : in std_logic;
slowed_clk : out std_logic);
end component;

component freq_div_20 
Port ( clk : in std_logic;
slowed_clk : out std_logic);
end component;

component shift_4
Port ( btn : in std_logic;
slowed_clk : in std_logic;
deb_out : out std_logic);
end component ;


begin

sq(hpos,vpos,refx,refy,assign_sq);

w1 : winning port map(reset,hpos,vpos,assign_sq,win_res,win);
f0 : freq_div_2 port map(vclk,ssclk);
f1 : freq_div_20 port map(vclk,slow);
d0 : shift_4 port map (VL,slow,dir(3));
d1 : shift_4 port map (VU,slow,dir(2));
d2 : shift_4 port map (VD,slow,dir(1));
d3 : shift_4 port map (VR,slow,dir(0));
m1 : mapp port map (hpos,vpos,win,assign_mapwin,assign_maze);


process(ssclk,reset,dir) 
--variable rgb : STD_LOGIC_VECTOR(7 downto 0);
begin
--
--   rgb:=rgb+"00000001";
--	if rgb="11111111" then
--	rgb:="00000000";
--   end if;
	
 if(reset='1') then
		refx<=16;
		refy<=16;
		hpos<=0;
		vpos<=0;
		vgahs<='0';
		vgavs<='0';
		vgar<="000";
		vgag<="000";
		vgab<="00";
elsif (ssclk'event and ssclk ='1') then

	                rgb:=rgb+"00000001";
						 if rgb="11111111" then
						 rgb:="00000000";
						 end if;
						 
	if(assign_sq='1') then
	if win='1' then
	vgar<="000";
	vgag<="000";
	vgab<="00";
	
	elsif dir(3)='1' then
         
						  vgar <= rgb(7 downto 5);
						  vgag <= rgb(4 downto 2);
						  vgab <= rgb(1 downto 0);
						
   elsif dir(2)='1' then
          
						  vgar <= rgb(7 downto 5);
						  vgag <= rgb(4 downto 2);
						  vgab <= rgb(1 downto 0);
						  
   elsif dir(1)='1' then
          
						  vgar <= rgb(7 downto 5);
						  vgag <= rgb(4 downto 2);
						  vgab <= rgb(1 downto 0);
						 
   elsif dir(0)='1' then
           
						  vgar <= rgb(7 downto 5);
						  vgag <= rgb(4 downto 2);
						  vgab <= rgb(1 downto 0);
					
			  else
					  vgar <= rgb(7 downto 5);
					  vgag <= rgb(4 downto 2);
					  vgab <= rgb(1 downto 0);
           end if;

	end if;
	if(assign_maze='1') then 
	vgar<="000";
	vgag<="000";
	vgab<="11";
	end if;
	if(assign_mapwin='1') then 
	--refx<=0;
	--refy<=0;
	--reset<=1;
	vgar<="000";
	vgag<="111";
	vgab<="00";
	end if;
	if(assign_sq='1' and assign_maze='1') then 
	refx<=16;
	refy<=16;
	end if;
--	if(assign_sq='1' and win_res='1') then 
--	refx<=16;
--	refy<=16;
--	end if;
	if(assign_sq='0' and assign_maze='0' and assign_mapwin='0')  then  
	vgar<="000";
	vgag<="000";
	vgab<="00";
   end if;
   --end if;
	if hpos < h_period  then
			hpos <= hpos+1;
		else 
			hpos<=0;
			if vpos < v_period  then
				vpos <= vpos+1;
	      else 
				vpos <= 0;
				if (dir(3)='1') then
				  refx <= refx-5;
--					if assign_sq='1' then
--						rgb:=rgb+"00000001";
--						if rgb="11111111" then
--						rgb:="00000000";
--						end if;
--					vgar <= rgb(7 downto 5);
--					vgag <= rgb(4 downto 2);
--					vgab <= rgb(1 downto 0);
--					end if;
				  elsif(dir(2)='1') then
				  refy <= refy-5;
--					if assign_sq='1' then
--						rgb:=rgb+"00000001";
--						if rgb="11111111" then
--						rgb:="00000000";
--						end if;
--					vgar <= rgb(7 downto 5);
--					vgag <= rgb(4 downto 2);
--					vgab <= rgb(1 downto 0);
--					end if;
				  elsif (dir(1)='1') then
				  refy <= refy+5;
--					if assign_sq='1' then
--						rgb:=rgb+"00000001";
--						if rgb="11111111" then
--						rgb:="00000000";
--						end if;
--					vgar <= rgb(7 downto 5);
--					vgag <= rgb(4 downto 2);
--					vgab <= rgb(1 downto 0);
--					end if;
				  elsif (dir(0)='1') then
				  refx <= refx+5;
--				  	if assign_sq='1' then
--						rgb:=rgb+"00000001";
--						if rgb="11111111" then
--						rgb:="00000000";
--						end if;
--					vgar <= rgb(7 downto 5);
--					vgag <= rgb(4 downto 2);
--					vgab <= rgb(1 downto 0);
--					end if;
				  else 
				  refx<=refx;
				  refy<=refy;
				  end if;
	      end if;
		end if;
	end if;
	
 IF((HPOS>H_DISP) OR (VPOS>V_DISP))THEN
	vgar<="000";
	vgag<="000";
	vgab<="00";
	END IF;
	
   if(hpos < H_DISP + H_FP OR hpos>= H_DISP + H_FP + H_PW) then
				vgahs <='1';
         else
				vgahs <= '0';
         end if;
            
         if(vpos < V_DISP + V_FP OR vpos >= V_DISP + V_FP + V_PW) then
				vgavs<= '1';
         else
				vgavs <= '0';
         end if;
	
end process;

end Behavioral;
